library verilog;
use verilog.vl_types.all;
entity NLC_1ch_1 is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        srdyi           : in     vl_logic;
        x_lin           : out    vl_logic_vector(20 downto 0);
        srdyo           : out    vl_logic;
        x_adc           : in     vl_logic_vector(20 downto 0);
        section_limit   : in     vl_logic_vector(19 downto 0);
        recip_stdev_4   : in     vl_logic_vector(31 downto 0);
        recip_stdev_3   : in     vl_logic_vector(31 downto 0);
        recip_stdev_2   : in     vl_logic_vector(31 downto 0);
        recip_stdev_1   : in     vl_logic_vector(31 downto 0);
        neg_mean_4      : in     vl_logic_vector(31 downto 0);
        neg_mean_3      : in     vl_logic_vector(31 downto 0);
        neg_mean_2      : in     vl_logic_vector(31 downto 0);
        neg_mean_1      : in     vl_logic_vector(31 downto 0);
        coeff_4_10      : in     vl_logic_vector(31 downto 0);
        coeff_4_9       : in     vl_logic_vector(31 downto 0);
        coeff_4_8       : in     vl_logic_vector(31 downto 0);
        coeff_4_7       : in     vl_logic_vector(31 downto 0);
        coeff_4_6       : in     vl_logic_vector(31 downto 0);
        coeff_4_5       : in     vl_logic_vector(31 downto 0);
        coeff_4_4       : in     vl_logic_vector(31 downto 0);
        coeff_4_3       : in     vl_logic_vector(31 downto 0);
        coeff_4_2       : in     vl_logic_vector(31 downto 0);
        coeff_4_1       : in     vl_logic_vector(31 downto 0);
        coeff_4_0       : in     vl_logic_vector(31 downto 0);
        coeff_3_10      : in     vl_logic_vector(31 downto 0);
        coeff_3_9       : in     vl_logic_vector(31 downto 0);
        coeff_3_8       : in     vl_logic_vector(31 downto 0);
        coeff_3_7       : in     vl_logic_vector(31 downto 0);
        coeff_3_6       : in     vl_logic_vector(31 downto 0);
        coeff_3_5       : in     vl_logic_vector(31 downto 0);
        coeff_3_4       : in     vl_logic_vector(31 downto 0);
        coeff_3_3       : in     vl_logic_vector(31 downto 0);
        coeff_3_2       : in     vl_logic_vector(31 downto 0);
        coeff_3_1       : in     vl_logic_vector(31 downto 0);
        coeff_3_0       : in     vl_logic_vector(31 downto 0);
        coeff_2_10      : in     vl_logic_vector(31 downto 0);
        coeff_2_9       : in     vl_logic_vector(31 downto 0);
        coeff_2_8       : in     vl_logic_vector(31 downto 0);
        coeff_2_7       : in     vl_logic_vector(31 downto 0);
        coeff_2_6       : in     vl_logic_vector(31 downto 0);
        coeff_2_5       : in     vl_logic_vector(31 downto 0);
        coeff_2_4       : in     vl_logic_vector(31 downto 0);
        coeff_2_3       : in     vl_logic_vector(31 downto 0);
        coeff_2_2       : in     vl_logic_vector(31 downto 0);
        coeff_2_1       : in     vl_logic_vector(31 downto 0);
        coeff_2_0       : in     vl_logic_vector(31 downto 0);
        coeff_1_10      : in     vl_logic_vector(31 downto 0);
        coeff_1_9       : in     vl_logic_vector(31 downto 0);
        coeff_1_8       : in     vl_logic_vector(31 downto 0);
        coeff_1_7       : in     vl_logic_vector(31 downto 0);
        coeff_1_6       : in     vl_logic_vector(31 downto 0);
        coeff_1_5       : in     vl_logic_vector(31 downto 0);
        coeff_1_4       : in     vl_logic_vector(31 downto 0);
        coeff_1_3       : in     vl_logic_vector(31 downto 0);
        coeff_1_2       : in     vl_logic_vector(31 downto 0);
        coeff_1_1       : in     vl_logic_vector(31 downto 0);
        coeff_1_0       : in     vl_logic_vector(31 downto 0)
    );
end NLC_1ch_1;
