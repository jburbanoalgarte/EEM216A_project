library verilog;
use verilog.vl_types.all;
entity NLC_4sec_10th_order_32ch_v0 is
    port(
        clk             : in     vl_logic;
        GlobalReset     : in     vl_logic;
        srdyo           : out    vl_logic;
        srdyi           : in     vl_logic;
        ch31_x_lin      : out    vl_logic_vector(20 downto 0);
        ch31_x_adc      : in     vl_logic_vector(20 downto 0);
        ch31_section_limit: in     vl_logic_vector(19 downto 0);
        ch31_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch31_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch30_x_lin      : out    vl_logic_vector(20 downto 0);
        ch30_x_adc      : in     vl_logic_vector(20 downto 0);
        ch30_section_limit: in     vl_logic_vector(19 downto 0);
        ch30_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch30_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch29_x_lin      : out    vl_logic_vector(20 downto 0);
        ch29_x_adc      : in     vl_logic_vector(20 downto 0);
        ch29_section_limit: in     vl_logic_vector(19 downto 0);
        ch29_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch29_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch28_x_lin      : out    vl_logic_vector(20 downto 0);
        ch28_x_adc      : in     vl_logic_vector(20 downto 0);
        ch28_section_limit: in     vl_logic_vector(19 downto 0);
        ch28_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch28_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch27_x_lin      : out    vl_logic_vector(20 downto 0);
        ch27_x_adc      : in     vl_logic_vector(20 downto 0);
        ch27_section_limit: in     vl_logic_vector(19 downto 0);
        ch27_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch27_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch26_x_lin      : out    vl_logic_vector(20 downto 0);
        ch26_x_adc      : in     vl_logic_vector(20 downto 0);
        ch26_section_limit: in     vl_logic_vector(19 downto 0);
        ch26_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch26_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch25_x_lin      : out    vl_logic_vector(20 downto 0);
        ch25_x_adc      : in     vl_logic_vector(20 downto 0);
        ch25_section_limit: in     vl_logic_vector(19 downto 0);
        ch25_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch25_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch24_x_lin      : out    vl_logic_vector(20 downto 0);
        ch24_x_adc      : in     vl_logic_vector(20 downto 0);
        ch24_section_limit: in     vl_logic_vector(19 downto 0);
        ch24_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch24_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch23_x_lin      : out    vl_logic_vector(20 downto 0);
        ch23_x_adc      : in     vl_logic_vector(20 downto 0);
        ch23_section_limit: in     vl_logic_vector(19 downto 0);
        ch23_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch23_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch22_x_lin      : out    vl_logic_vector(20 downto 0);
        ch22_x_adc      : in     vl_logic_vector(20 downto 0);
        ch22_section_limit: in     vl_logic_vector(19 downto 0);
        ch22_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch22_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch21_x_lin      : out    vl_logic_vector(20 downto 0);
        ch21_x_adc      : in     vl_logic_vector(20 downto 0);
        ch21_section_limit: in     vl_logic_vector(19 downto 0);
        ch21_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch21_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch20_x_lin      : out    vl_logic_vector(20 downto 0);
        ch20_x_adc      : in     vl_logic_vector(20 downto 0);
        ch20_section_limit: in     vl_logic_vector(19 downto 0);
        ch20_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch20_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch19_x_lin      : out    vl_logic_vector(20 downto 0);
        ch19_x_adc      : in     vl_logic_vector(20 downto 0);
        ch19_section_limit: in     vl_logic_vector(19 downto 0);
        ch19_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch19_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch18_x_lin      : out    vl_logic_vector(20 downto 0);
        ch18_x_adc      : in     vl_logic_vector(20 downto 0);
        ch18_section_limit: in     vl_logic_vector(19 downto 0);
        ch18_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch18_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch17_x_lin      : out    vl_logic_vector(20 downto 0);
        ch17_x_adc      : in     vl_logic_vector(20 downto 0);
        ch17_section_limit: in     vl_logic_vector(19 downto 0);
        ch17_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch17_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch16_x_lin      : out    vl_logic_vector(20 downto 0);
        ch16_x_adc      : in     vl_logic_vector(20 downto 0);
        ch16_section_limit: in     vl_logic_vector(19 downto 0);
        ch16_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch16_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch15_x_lin      : out    vl_logic_vector(20 downto 0);
        ch15_x_adc      : in     vl_logic_vector(20 downto 0);
        ch15_section_limit: in     vl_logic_vector(19 downto 0);
        ch15_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch15_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch14_x_lin      : out    vl_logic_vector(20 downto 0);
        ch14_x_adc      : in     vl_logic_vector(20 downto 0);
        ch14_section_limit: in     vl_logic_vector(19 downto 0);
        ch14_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch14_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch13_x_lin      : out    vl_logic_vector(20 downto 0);
        ch13_x_adc      : in     vl_logic_vector(20 downto 0);
        ch13_section_limit: in     vl_logic_vector(19 downto 0);
        ch13_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch13_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch12_x_lin      : out    vl_logic_vector(20 downto 0);
        ch12_x_adc      : in     vl_logic_vector(20 downto 0);
        ch12_section_limit: in     vl_logic_vector(19 downto 0);
        ch12_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch12_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch11_x_lin      : out    vl_logic_vector(20 downto 0);
        ch11_x_adc      : in     vl_logic_vector(20 downto 0);
        ch11_section_limit: in     vl_logic_vector(19 downto 0);
        ch11_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch11_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch10_x_lin      : out    vl_logic_vector(20 downto 0);
        ch10_x_adc      : in     vl_logic_vector(20 downto 0);
        ch10_section_limit: in     vl_logic_vector(19 downto 0);
        ch10_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch10_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch9_x_lin       : out    vl_logic_vector(20 downto 0);
        ch9_x_adc       : in     vl_logic_vector(20 downto 0);
        ch9_section_limit: in     vl_logic_vector(19 downto 0);
        ch9_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch9_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch8_x_lin       : out    vl_logic_vector(20 downto 0);
        ch8_x_adc       : in     vl_logic_vector(20 downto 0);
        ch8_section_limit: in     vl_logic_vector(19 downto 0);
        ch8_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch8_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch7_x_lin       : out    vl_logic_vector(20 downto 0);
        ch7_x_adc       : in     vl_logic_vector(20 downto 0);
        ch7_section_limit: in     vl_logic_vector(19 downto 0);
        ch7_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch7_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch6_x_lin       : out    vl_logic_vector(20 downto 0);
        ch6_x_adc       : in     vl_logic_vector(20 downto 0);
        ch6_section_limit: in     vl_logic_vector(19 downto 0);
        ch6_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch6_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch5_x_lin       : out    vl_logic_vector(20 downto 0);
        ch5_x_adc       : in     vl_logic_vector(20 downto 0);
        ch5_section_limit: in     vl_logic_vector(19 downto 0);
        ch5_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch5_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch4_x_lin       : out    vl_logic_vector(20 downto 0);
        ch4_x_adc       : in     vl_logic_vector(20 downto 0);
        ch4_section_limit: in     vl_logic_vector(19 downto 0);
        ch4_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch4_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch3_x_lin       : out    vl_logic_vector(20 downto 0);
        ch3_x_adc       : in     vl_logic_vector(20 downto 0);
        ch3_section_limit: in     vl_logic_vector(19 downto 0);
        ch3_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch3_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch2_x_lin       : out    vl_logic_vector(20 downto 0);
        ch2_x_adc       : in     vl_logic_vector(20 downto 0);
        ch2_section_limit: in     vl_logic_vector(19 downto 0);
        ch2_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch2_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch1_x_lin       : out    vl_logic_vector(20 downto 0);
        ch1_x_adc       : in     vl_logic_vector(20 downto 0);
        ch1_section_limit: in     vl_logic_vector(19 downto 0);
        ch1_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch1_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0);
        ch0_x_lin       : out    vl_logic_vector(20 downto 0);
        ch0_x_adc       : in     vl_logic_vector(20 downto 0);
        ch0_section_limit: in     vl_logic_vector(19 downto 0);
        ch0_select_section_coefficients_stdev_4_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_stdev_3_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_stdev_2_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_stdev_1_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_mean_4_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_mean_3_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_mean_2_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_mean_1_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_9_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_8_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_7_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_6_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_5_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_4_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_3_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_2_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_10_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_1_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_4_0_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_9_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_8_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_7_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_6_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_5_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_4_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_3_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_2_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_10_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_1_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_3_0_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_9_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_8_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_7_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_6_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_5_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_4_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_3_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_2_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_10_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_1_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_2_0_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_9_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_8_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_7_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_6_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_5_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_4_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_3_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_2_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_10_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_1_porty: in     vl_logic_vector(31 downto 0);
        ch0_select_section_coefficients_coeff_1_0_porty: in     vl_logic_vector(31 downto 0)
    );
end NLC_4sec_10th_order_32ch_v0;
