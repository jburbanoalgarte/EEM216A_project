library verilog;
use verilog.vl_types.all;
entity comparator is
    port(
        clk             : in     vl_logic;
        GlobalReset     : in     vl_logic;
        x_adc_latched   : in     vl_logic_vector(20 downto 0);
        section_limit   : in     vl_logic_vector(19 downto 0);
        coeff1_0        : in     vl_logic_vector(31 downto 0);
        coeff1_1        : in     vl_logic_vector(31 downto 0);
        coeff1_2        : in     vl_logic_vector(31 downto 0);
        coeff1_3        : in     vl_logic_vector(31 downto 0);
        coeff1_4        : in     vl_logic_vector(31 downto 0);
        coeff1_5        : in     vl_logic_vector(31 downto 0);
        coeff1_6        : in     vl_logic_vector(31 downto 0);
        coeff1_7        : in     vl_logic_vector(31 downto 0);
        coeff1_8        : in     vl_logic_vector(31 downto 0);
        coeff1_9        : in     vl_logic_vector(31 downto 0);
        coeff1_10       : in     vl_logic_vector(31 downto 0);
        mean1           : in     vl_logic_vector(31 downto 0);
        std1            : in     vl_logic_vector(31 downto 0);
        coeff2_0        : in     vl_logic_vector(31 downto 0);
        coeff2_1        : in     vl_logic_vector(31 downto 0);
        coeff2_2        : in     vl_logic_vector(31 downto 0);
        coeff2_3        : in     vl_logic_vector(31 downto 0);
        coeff2_4        : in     vl_logic_vector(31 downto 0);
        coeff2_5        : in     vl_logic_vector(31 downto 0);
        coeff2_6        : in     vl_logic_vector(31 downto 0);
        coeff2_7        : in     vl_logic_vector(31 downto 0);
        coeff2_8        : in     vl_logic_vector(31 downto 0);
        coeff2_9        : in     vl_logic_vector(31 downto 0);
        coeff2_10       : in     vl_logic_vector(31 downto 0);
        mean2           : in     vl_logic_vector(31 downto 0);
        std2            : in     vl_logic_vector(31 downto 0);
        coeff3_0        : in     vl_logic_vector(31 downto 0);
        coeff3_1        : in     vl_logic_vector(31 downto 0);
        coeff3_2        : in     vl_logic_vector(31 downto 0);
        coeff3_3        : in     vl_logic_vector(31 downto 0);
        coeff3_4        : in     vl_logic_vector(31 downto 0);
        coeff3_5        : in     vl_logic_vector(31 downto 0);
        coeff3_6        : in     vl_logic_vector(31 downto 0);
        coeff3_7        : in     vl_logic_vector(31 downto 0);
        coeff3_8        : in     vl_logic_vector(31 downto 0);
        coeff3_9        : in     vl_logic_vector(31 downto 0);
        coeff3_10       : in     vl_logic_vector(31 downto 0);
        mean3           : in     vl_logic_vector(31 downto 0);
        std3            : in     vl_logic_vector(31 downto 0);
        coeff4_0        : in     vl_logic_vector(31 downto 0);
        coeff4_1        : in     vl_logic_vector(31 downto 0);
        coeff4_2        : in     vl_logic_vector(31 downto 0);
        coeff4_3        : in     vl_logic_vector(31 downto 0);
        coeff4_4        : in     vl_logic_vector(31 downto 0);
        coeff4_5        : in     vl_logic_vector(31 downto 0);
        coeff4_6        : in     vl_logic_vector(31 downto 0);
        coeff4_7        : in     vl_logic_vector(31 downto 0);
        coeff4_8        : in     vl_logic_vector(31 downto 0);
        coeff4_9        : in     vl_logic_vector(31 downto 0);
        coeff4_10       : in     vl_logic_vector(31 downto 0);
        mean4           : in     vl_logic_vector(31 downto 0);
        std4            : in     vl_logic_vector(31 downto 0);
        coeff0          : out    vl_logic_vector(31 downto 0);
        coeff1          : out    vl_logic_vector(31 downto 0);
        coeff2          : out    vl_logic_vector(31 downto 0);
        coeff3          : out    vl_logic_vector(31 downto 0);
        coeff4          : out    vl_logic_vector(31 downto 0);
        coeff5          : out    vl_logic_vector(31 downto 0);
        coeff6          : out    vl_logic_vector(31 downto 0);
        coeff7          : out    vl_logic_vector(31 downto 0);
        coeff8          : out    vl_logic_vector(31 downto 0);
        coeff9          : out    vl_logic_vector(31 downto 0);
        coeff10         : out    vl_logic_vector(31 downto 0);
        mean            : out    vl_logic_vector(31 downto 0);
        std             : out    vl_logic_vector(31 downto 0)
    );
end comparator;
