library verilog;
use verilog.vl_types.all;
entity test_NLC_4sec_10th_order_32ch_v0 is
end test_NLC_4sec_10th_order_32ch_v0;
