library verilog;
use verilog.vl_types.all;
entity NLC_1ch is
    port(
        clk             : in     vl_logic;
        reset           : in     vl_logic;
        srdyi           : in     vl_logic;
        srdyo           : out    vl_logic;
        ch31_x_adc      : in     vl_logic_vector(20 downto 0);
        ch31_x_lin      : out    vl_logic_vector(20 downto 0);
        ch31_section_limit: in     vl_logic_vector(19 downto 0);
        ch31_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch31_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch31_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch31_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch31_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch31_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch31_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch31_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch31_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch30_x_adc      : in     vl_logic_vector(20 downto 0);
        ch30_x_lin      : out    vl_logic_vector(20 downto 0);
        ch30_section_limit: in     vl_logic_vector(19 downto 0);
        ch30_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch30_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch30_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch30_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch30_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch30_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch30_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch30_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch30_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch29_x_adc      : in     vl_logic_vector(20 downto 0);
        ch29_x_lin      : out    vl_logic_vector(20 downto 0);
        ch29_section_limit: in     vl_logic_vector(19 downto 0);
        ch29_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch29_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch29_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch29_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch29_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch29_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch29_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch29_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch29_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch28_x_adc      : in     vl_logic_vector(20 downto 0);
        ch28_x_lin      : out    vl_logic_vector(20 downto 0);
        ch28_section_limit: in     vl_logic_vector(19 downto 0);
        ch28_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch28_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch28_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch28_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch28_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch28_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch28_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch28_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch28_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch27_x_adc      : in     vl_logic_vector(20 downto 0);
        ch27_x_lin      : out    vl_logic_vector(20 downto 0);
        ch27_section_limit: in     vl_logic_vector(19 downto 0);
        ch27_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch27_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch27_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch27_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch27_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch27_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch27_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch27_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch27_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch26_x_adc      : in     vl_logic_vector(20 downto 0);
        ch26_x_lin      : out    vl_logic_vector(20 downto 0);
        ch26_section_limit: in     vl_logic_vector(19 downto 0);
        ch26_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch26_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch26_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch26_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch26_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch26_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch26_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch26_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch26_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch25_x_adc      : in     vl_logic_vector(20 downto 0);
        ch25_x_lin      : out    vl_logic_vector(20 downto 0);
        ch25_section_limit: in     vl_logic_vector(19 downto 0);
        ch25_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch25_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch25_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch25_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch25_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch25_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch25_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch25_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch25_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch24_x_adc      : in     vl_logic_vector(20 downto 0);
        ch24_x_lin      : out    vl_logic_vector(20 downto 0);
        ch24_section_limit: in     vl_logic_vector(19 downto 0);
        ch24_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch24_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch24_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch24_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch24_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch24_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch24_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch24_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch24_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch23_x_adc      : in     vl_logic_vector(20 downto 0);
        ch23_x_lin      : out    vl_logic_vector(20 downto 0);
        ch23_section_limit: in     vl_logic_vector(19 downto 0);
        ch23_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch23_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch23_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch23_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch23_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch23_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch23_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch23_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch23_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch22_x_adc      : in     vl_logic_vector(20 downto 0);
        ch22_x_lin      : out    vl_logic_vector(20 downto 0);
        ch22_section_limit: in     vl_logic_vector(19 downto 0);
        ch22_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch22_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch22_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch22_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch22_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch22_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch22_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch22_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch22_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch21_x_adc      : in     vl_logic_vector(20 downto 0);
        ch21_x_lin      : out    vl_logic_vector(20 downto 0);
        ch21_section_limit: in     vl_logic_vector(19 downto 0);
        ch21_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch21_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch21_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch21_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch21_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch21_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch21_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch21_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch21_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch20_x_adc      : in     vl_logic_vector(20 downto 0);
        ch20_x_lin      : out    vl_logic_vector(20 downto 0);
        ch20_section_limit: in     vl_logic_vector(19 downto 0);
        ch20_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch20_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch20_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch20_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch20_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch20_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch20_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch20_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch20_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch19_x_adc      : in     vl_logic_vector(20 downto 0);
        ch19_x_lin      : out    vl_logic_vector(20 downto 0);
        ch19_section_limit: in     vl_logic_vector(19 downto 0);
        ch19_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch19_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch19_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch19_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch19_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch19_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch19_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch19_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch19_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch18_x_adc      : in     vl_logic_vector(20 downto 0);
        ch18_x_lin      : out    vl_logic_vector(20 downto 0);
        ch18_section_limit: in     vl_logic_vector(19 downto 0);
        ch18_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch18_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch18_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch18_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch18_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch18_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch18_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch18_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch18_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch17_x_adc      : in     vl_logic_vector(20 downto 0);
        ch17_x_lin      : out    vl_logic_vector(20 downto 0);
        ch17_section_limit: in     vl_logic_vector(19 downto 0);
        ch17_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch17_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch17_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch17_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch17_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch17_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch17_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch17_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch17_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch16_x_adc      : in     vl_logic_vector(20 downto 0);
        ch16_x_lin      : out    vl_logic_vector(20 downto 0);
        ch16_section_limit: in     vl_logic_vector(19 downto 0);
        ch16_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch16_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch16_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch16_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch16_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch16_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch16_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch16_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch16_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch15_x_adc      : in     vl_logic_vector(20 downto 0);
        ch15_x_lin      : out    vl_logic_vector(20 downto 0);
        ch15_section_limit: in     vl_logic_vector(19 downto 0);
        ch15_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch15_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch15_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch15_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch15_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch15_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch15_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch15_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch15_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch14_x_adc      : in     vl_logic_vector(20 downto 0);
        ch14_x_lin      : out    vl_logic_vector(20 downto 0);
        ch14_section_limit: in     vl_logic_vector(19 downto 0);
        ch14_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch14_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch14_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch14_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch14_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch14_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch14_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch14_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch14_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch13_x_adc      : in     vl_logic_vector(20 downto 0);
        ch13_x_lin      : out    vl_logic_vector(20 downto 0);
        ch13_section_limit: in     vl_logic_vector(19 downto 0);
        ch13_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch13_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch13_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch13_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch13_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch13_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch13_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch13_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch13_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch12_x_adc      : in     vl_logic_vector(20 downto 0);
        ch12_x_lin      : out    vl_logic_vector(20 downto 0);
        ch12_section_limit: in     vl_logic_vector(19 downto 0);
        ch12_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch12_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch12_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch12_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch12_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch12_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch12_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch12_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch12_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch11_x_adc      : in     vl_logic_vector(20 downto 0);
        ch11_x_lin      : out    vl_logic_vector(20 downto 0);
        ch11_section_limit: in     vl_logic_vector(19 downto 0);
        ch11_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch11_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch11_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch11_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch11_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch11_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch11_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch11_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch11_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch10_x_adc      : in     vl_logic_vector(20 downto 0);
        ch10_x_lin      : out    vl_logic_vector(20 downto 0);
        ch10_section_limit: in     vl_logic_vector(19 downto 0);
        ch10_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch10_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch10_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch10_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch10_neg_mean_4 : in     vl_logic_vector(31 downto 0);
        ch10_neg_mean_3 : in     vl_logic_vector(31 downto 0);
        ch10_neg_mean_2 : in     vl_logic_vector(31 downto 0);
        ch10_neg_mean_1 : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_10 : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_9  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_8  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_7  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_6  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_5  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_4  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_3  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_2  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_1  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_4_0  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_10 : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_9  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_8  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_7  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_6  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_5  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_4  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_3  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_2  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_1  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_3_0  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_10 : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_9  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_8  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_7  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_6  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_5  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_4  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_3  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_2  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_1  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_2_0  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_10 : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_9  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_8  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_7  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_6  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_5  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_4  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_3  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_2  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_1  : in     vl_logic_vector(31 downto 0);
        ch10_coeff_1_0  : in     vl_logic_vector(31 downto 0);
        ch9_x_adc       : in     vl_logic_vector(20 downto 0);
        ch9_x_lin       : out    vl_logic_vector(20 downto 0);
        ch9_section_limit: in     vl_logic_vector(19 downto 0);
        ch9_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch9_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch9_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch9_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch9_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch9_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch9_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch9_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch9_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch8_x_adc       : in     vl_logic_vector(20 downto 0);
        ch8_x_lin       : out    vl_logic_vector(20 downto 0);
        ch8_section_limit: in     vl_logic_vector(19 downto 0);
        ch8_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch8_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch8_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch8_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch8_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch8_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch8_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch8_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch8_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch7_x_adc       : in     vl_logic_vector(20 downto 0);
        ch7_x_lin       : out    vl_logic_vector(20 downto 0);
        ch7_section_limit: in     vl_logic_vector(19 downto 0);
        ch7_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch7_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch7_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch7_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch7_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch7_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch7_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch7_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch7_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch6_x_adc       : in     vl_logic_vector(20 downto 0);
        ch6_x_lin       : out    vl_logic_vector(20 downto 0);
        ch6_section_limit: in     vl_logic_vector(19 downto 0);
        ch6_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch6_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch6_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch6_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch6_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch6_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch6_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch6_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch6_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch5_x_adc       : in     vl_logic_vector(20 downto 0);
        ch5_x_lin       : out    vl_logic_vector(20 downto 0);
        ch5_section_limit: in     vl_logic_vector(19 downto 0);
        ch5_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch5_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch5_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch5_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch5_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch5_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch5_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch5_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch5_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch4_x_adc       : in     vl_logic_vector(20 downto 0);
        ch4_x_lin       : out    vl_logic_vector(20 downto 0);
        ch4_section_limit: in     vl_logic_vector(19 downto 0);
        ch4_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch4_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch4_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch4_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch4_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch4_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch4_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch4_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch4_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch3_x_adc       : in     vl_logic_vector(20 downto 0);
        ch3_x_lin       : out    vl_logic_vector(20 downto 0);
        ch3_section_limit: in     vl_logic_vector(19 downto 0);
        ch3_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch3_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch3_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch3_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch3_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch3_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch3_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch3_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch3_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch2_x_adc       : in     vl_logic_vector(20 downto 0);
        ch2_x_lin       : out    vl_logic_vector(20 downto 0);
        ch2_section_limit: in     vl_logic_vector(19 downto 0);
        ch2_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch2_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch2_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch2_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch2_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch2_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch2_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch2_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch2_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch1_x_adc       : in     vl_logic_vector(20 downto 0);
        ch1_x_lin       : out    vl_logic_vector(20 downto 0);
        ch1_section_limit: in     vl_logic_vector(19 downto 0);
        ch1_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch1_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch1_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch1_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch1_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch1_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch1_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch1_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch1_coeff_1_0   : in     vl_logic_vector(31 downto 0);
        ch0_x_adc       : in     vl_logic_vector(20 downto 0);
        ch0_x_lin       : out    vl_logic_vector(20 downto 0);
        ch0_section_limit: in     vl_logic_vector(19 downto 0);
        ch0_recip_stdev_4: in     vl_logic_vector(31 downto 0);
        ch0_recip_stdev_3: in     vl_logic_vector(31 downto 0);
        ch0_recip_stdev_2: in     vl_logic_vector(31 downto 0);
        ch0_recip_stdev_1: in     vl_logic_vector(31 downto 0);
        ch0_neg_mean_4  : in     vl_logic_vector(31 downto 0);
        ch0_neg_mean_3  : in     vl_logic_vector(31 downto 0);
        ch0_neg_mean_2  : in     vl_logic_vector(31 downto 0);
        ch0_neg_mean_1  : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_10  : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_9   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_8   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_7   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_6   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_5   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_4   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_3   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_2   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_1   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_4_0   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_10  : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_9   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_8   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_7   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_6   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_5   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_4   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_3   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_2   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_1   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_3_0   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_10  : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_9   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_8   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_7   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_6   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_5   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_4   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_3   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_2   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_1   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_2_0   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_10  : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_9   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_8   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_7   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_6   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_5   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_4   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_3   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_2   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_1   : in     vl_logic_vector(31 downto 0);
        ch0_coeff_1_0   : in     vl_logic_vector(31 downto 0)
    );
end NLC_1ch;
